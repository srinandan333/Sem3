//program for 16-bit barrel shifter(only right shift)
module mux2_1(input wire x,y,s, output wire z);
    assign z = (s==0)?x:y;
endmodule

module barrelshifter(input wire [15:0] i, input wire [3:0] s, output wire [15:0] o);
    wire [15:0] c0, c1, c2;
    mux2_1 a0(i[15],1'b0,s[3],c0[15]);
    mux2_1 a1(i[14],1'b0,s[3],c0[14]);
    mux2_1 a2(i[13],1'b0,s[3],c0[13]);
    mux2_1 a3(i[12],1'b0,s[3],c0[12]);
    mux2_1 a4(i[11],1'b0,s[3],c0[11]);
    mux2_1 a5(i[10],1'b0,s[3],c0[10]);
    mux2_1 a6(i[9],1'b0,s[3],c0[9]);
    mux2_1 a7(i[8],1'b0,s[3],c0[8]);
    mux2_1 a8(i[7],i[15],s[3],c0[7]);
    mux2_1 a9(i[6],i[14],s[3],c0[6]);
    mux2_1 a10(i[5],i[13],s[3],c0[5]);
    mux2_1 a11(i[4],i[12],s[3],c0[4]);
    mux2_1 a12(i[3],i[11],s[3],c0[3]);
    mux2_1 a13(i[2],i[10],s[3],c0[2]);
    mux2_1 a14(i[1],i[9],s[3],c0[1]);
    mux2_1 a15(i[0],i[8],s[3],c0[0]);

    mux2_1 b0(c0[15],1'b0,s[2],c1[15]);
    mux2_1 b1(c0[14],1'b0,s[2],c1[14]);
    mux2_1 b2(c0[13],1'b0,s[2],c1[13]);
    mux2_1 b3(c0[12],1'b0,s[2],c1[12]);
    mux2_1 b4(c0[11],c0[15],s[2],c1[11]);
    mux2_1 b5(c0[10],c0[14],s[2],c1[10]);
    mux2_1 b6(c0[9],c0[13],s[2],c1[9]);
    mux2_1 b7(c0[8],c0[12],s[2],c1[8]);
    mux2_1 b8(c0[7],c0[11],s[2],c1[7]);
    mux2_1 b9(c0[6],c0[10],s[2],c1[6]);
    mux2_1 b10(c0[5],c0[9],s[2],c1[5]);
    mux2_1 b11(c0[4],c0[8],s[2],c1[4]);
    mux2_1 b12(c0[3],c0[7],s[2],c1[3]);
    mux2_1 b13(c0[2],c0[6],s[2],c1[2]);
    mux2_1 b14(c0[1],c0[5],s[2],c1[1]);
    mux2_1 b15(c0[0],c0[4],s[2],c1[0]);

    mux2_1 c0(c1[15],1'b0,s[1],c2[15]);
    mux2_1 c1(c1[14],1'b0,s[1],c2[14]);
    mux2_1 c2(c1[13],c1[15],s[1],c2[13]);
    mux2_1 c3(c1[12],c1[14],s[1],c2[12]);
    mux2_1 c4(c1[11],c1[13],s[1],c2[11]);
    mux2_1 c5(c1[10],c1[12],s[1],c2[10]);
    mux2_1 c6(c1[9],c1[11],s[1],c2[9]);
    mux2_1 c7(c1[8],c1[10],s[1],c2[8]);
    mux2_1 c8(c1[7],c1[9],s[1],c2[7]);
    mux2_1 c9(c1[6],c1[8],s[1],c2[6]);
    mux2_1 c10(c1[5],c1[7],s[1],c2[5]);
    mux2_1 c11(c1[4],c1[6],s[1],c2[4]);
    mux2_1 c12(c1[3],c1[5],s[1],c2[3]);
    mux2_1 c13(c1[2],c1[4],s[1],c2[2]);
    mux2_1 c14(c1[1],c1[3],s[1],c2[1]);
    mux2_1 c15(c1[0],c1[2],s[1],c2[0]);

    mux2_1 d0(c2[15],1'b0,s[0],o[15]);
    mux2_1 d1(c2[14],c2[15],s[0],o[14]);
    mux2_1 d2(c2[13],c2[14],s[0],o[13]);
    mux2_1 d3(c2[12],c2[13],s[0],o[12]);
    mux2_1 d4(c2[11],c2[12],s[0],o[11]);
    mux2_1 d5(c2[10],c2[11],s[0],o[10]);
    mux2_1 d6(c2[9],c2[10],s[0],o[9]);
    mux2_1 d7(c2[8],c2[9],s[0],o[8]);
    mux2_1 d8(c2[7],c2[8],s[0],o[7]);
    mux2_1 d9(c2[6],c2[7],s[0],o[6]);
    mux2_1 d10(c2[5],c2[6],s[0],o[5]);
    mux2_1 d11(c2[4],c2[5],s[0],o[4]);
    mux2_1 d12(c2[3],c2[4],s[0],o[3]);
    mux2_1 d13(c2[2],c2[3],s[0],o[2]);
    mux2_1 d14(c2[1],c2[2],s[0],o[1]);
    mux2_1 d15(c2[0],c2[1],s[0],o[0]);
endmodule



    